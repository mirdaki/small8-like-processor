-- Matthew Booe

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package eight_busses is    

   type eight_bus_input is array(NATURAL range <>) of std_logic_vector(7 downto 0);
	
end eight_busses;

package body eight_busses is
   -- subprogram bodies here
end eight_busses;